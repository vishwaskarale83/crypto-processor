`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/02/2020 04:03:49 PM
// Design Name: 
// Module Name: key_generator
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Key_generator(clk,rst,randomize,AES_key_new,private_key_new,AES_key_gen,private_key_gen,private_key,AES_key_final,N);
	
	parameter WIDTH = 256;
	parameter temp_size = 256;
	parameter public_key = 64'd65537;
	parameter R = 128'd11980692079448174547167670;
	    
	input rst,clk,randomize;
	input private_key_new;
    input AES_key_new;
	
	output reg [127:0] private_key;
	output reg [127:0] N;
    output reg private_key_gen; 

	output wire [127:0] AES_key_final;
	//output wire randomize_complete;
    output AES_key_gen;
       
    integer k;
    	
    reg [8:0] storage1;
    reg [4:0] storage3;
    reg [4:0] storage4;
    reg [255:0] storage;
    reg [127:0] var = 128'd244155625894036;
    reg [127:0] M,product;
    
    reg [15:0] p3 = 16'd55633;
    reg [15:0] p4 = 16'd35837;
        
    AES_key_generator AES_key(
        .clk(clk),
        .new(AES_key_new),
        .done(AES_key_gen),
        .randomizer(AES_key_final),
        .p1(p3),
        .p2(p4),
        .continue(randomize)
        //.randomize_complete(randomize_complete)
    );

always@(posedge clk) begin


    if(rst == 0 && randomize == 1) begin   
        storage1 = AES_key_final[12:4];
        
        storage3[4:0] = AES_key_final[113:109];
        
        if (storage3 == 31) 
            storage3 = storage3-1;
        
        storage4[4:0] = AES_key_final[123:119];
        
        if (storage4 == 31) 
            storage4 = storage4-1;
        
        if (storage3 == storage4) begin
            if(storage3 == 0)
                storage3 = storage3 + 1;
            else 
                storage3 = storage3 - 1;
        end
    end
    
    if (private_key_new == 1) begin
        private_key = 0;
        private_key_gen = 0;
        N = 0;
    end
    
    if (private_key_new == 0) begin
        private_key = storage[255:128];
        N = storage[127:0];
        private_key_gen = 1;
    end
end

always@(*) begin
    case(storage1)
        0 : storage = 256'h00811fc3302c98543757011355524861526f40ad9afe67f19acde65695cbd1dd;
        1 : storage = 256'h121af97e39cda196ac4078f6e703ae79135427dad0f2a61df4fccc56b486d923;
        2 : storage = 256'h06a80e748815568de2f7f64ad6016fc1075f9cfc07ba357f68964987448cf1b9;
        3 : storage = 256'h17dce7f8240f812aa23455c8273892094921813d53ecab68210ac49ed1d7870f;
        4 : storage = 256'h381a8dbcda8291a3355870504867ac5198c1e2da1e53a3eba02ec1fe860b90db;
        5 : storage = 256'h03008bee2c7fce6a0872306035c1c25935d4a3ce70e79ea2ab62c906f429f2b7;
        6 : storage = 256'h04a4eb17d043e79c33d1516294d3be610bf0928161207ef073aacfdbff82789b;
        7 : storage = 256'h117e43a455df08211532593ff4ca610114a57a46db9cd9e76da1f1aa2d45ffad;
        8 : storage = 256'h61712f61799db8153872bd75f36983c1837f7776bcf6f6988de70714dcc3d721;
        9 : storage = 256'h0b379c19021b0a33f958243fd67933c1129f9c7e6ce6b24a30f2a165d54ebffd;
        10 : storage = 256'h27deb6f076fa39e40de1ca00741e69e171aa8ca9f5dfab875f0cfc77d4d373a7;
        11 : storage = 256'h111daef262d51b7e957669cbc6e68e5971513b4d30a1be9182c45edd2f229a9f;
        12 : storage = 256'h00dbc77b1bb65ee1124de383f96b81410da4a54cec79d4444f08b9940aada341;
        13 : storage = 256'h1d324b6d3b6a9ca0f6b978455a50d8c125e004b336e3615048b21910b6a65bef;
        14 : storage = 256'h0ee51c5c9eda7e51c74bc9150785d7d11991d2666a8bd1dec96ac95ff1d624c9;
        15 : storage = 256'h2d1f8eadbf09df92173771be025fa1d17073872fe431bfe990e5ef77fd90185f;
        16 : storage = 256'h1062aec9cb22c46aba9dca57377c1f0160b7b2a1db71de0db430d54ae2cdfbe5;
        17 : storage = 256'h422282d29df878c43affbe1ae538d7115c26e92dc1d0d07870f53246be999807;
        18 : storage = 256'h05bf97933f1078bf9cbb14f93a742d990a2c8bc15ab23e19ab9b1efdab10eb9b;
        19 : storage = 256'h3bf72a6783047d6d49d1f1d64a28877168e7bac7c4ee31d9035eb07167ba7c87;
        20 : storage = 256'h270546567fe819614889a53d241aad0166d9eb3321ebd54528e2ce14165850c7;
        21 : storage = 256'h1dc0511dd8cbe0904b38056609892db1292e9cf1cfc1d9342437c81d66e085b3;
        22 : storage = 256'h1cd53ff849c52f6976f0ff8b02e658115e4e95bbab2f0b7fbe250c3ed3b6b689;
        23 : storage = 256'h3cd769761bdfee736b554d862bf16e01626b62376965dc76bb11191bff9bdb65;
        24 : storage = 256'h7f429925741b67bdac9fb7399c5ee6d184dc0130e59d4935078cf449b6fcdc61;
        25 : storage = 256'h0b09f8713b9e2f54ebe47f9b5491f2f96bd58c8120c157d9210ce1a6157212d3;
        26 : storage = 256'h00c68415d7bd101549700db548d02e710257bd35d8985f7a1c505b43668cc4c1;
        27 : storage = 256'h13c4512a1e645b579a773988942c17a95a5b9e0ce2506b1161665faff582fe27;
        28 : storage = 256'h4c4e64fd16a276e335d28ae4ff587b816fa81efa0dab6fffc068498271286d5d;
        29 : storage = 256'h44d1e3f1c35a687955e50faaf9dad0e185bd729773721b6c2f25a0062a042d6f;
        30 : storage = 256'h0b1ad903b7af731f96f5c359ca36ce9115a6d8c9fbfcd298956044ece4ac0e89;
        31 : storage = 256'h00811fc3302c98543757011355524861526f40ad9afe67f19acde65695cbd1dd;
        32 : storage = 256'h0fc47525f3531fbdb333f1637bf44f0110c0ddf9ecfa913d185253c298146b0f;
        33 : storage = 256'h00c2d3001a2af8d6bd12674d4da1928106641be9dcef6f327ff5ff80db8cfabd;
        34 : storage = 256'h2c2800c5b77cc50180cf51483bc2e3213f6310c0d9d99a749bf589b203c9d22b;
        35 : storage = 256'h061546a164f2d426653034353f2806f184677269388eee00173730535af320a7;
        36 : storage = 256'h1c9df7496f3019daeb9734af5408edc12ea884849d310bde5d17b981f6015973;
        37 : storage = 256'h056b6af8b956690804a7d01c1f1945510a59511e196dbf33ac97eba82ce1df67;
        38 : storage = 256'h023e412d8bbc948e1ca4df15db1f924111e53e99690d80a1beeec0c112f75b01;
        39 : storage = 256'h50bb68596a762eb1136709a1dd3386a171fa2bde6b6fa15e4477bbcbd1ff5ac5;
        40 : storage = 256'h039da2740844df6aa3a8a4b4140f0e01102460d94389d477903bd88193721691;
        41 : storage = 256'h26b05441fa797fb114f9814623e0f78162857af844b5b2489ab99e11d9e5cc23;
        42 : storage = 256'h4fedd9d326dfa2236f69a8fa655f9ff16238102bdb3ec173845ff52a276c55fb;
        43 : storage = 256'h0166207f2ce2dcdd9a9f7801aa37ec210bd349c68696b155187f56839aaa3b65;
        44 : storage = 256'h1c57c8eef87f7abad3a1748cf377922120d420c98aaa832abdb6a3641591368b;
        45 : storage = 256'h111080f4f29036718f3e9d5d54193f611629a95384a003bededde0953d588c0d;
        46 : storage = 256'h53e12b6aa2acc70fafd8bd0c07aeef016177e6330bcc7b28c9b0ad3fb200c2bb;
        47 : storage = 256'h29c33c4e740e0dd9df42519d9125760153d4bbea1457ed8fdad16bea338c7719;
        48 : storage = 256'h27c8ae73e29c4b00fca0795393f2b6d14fdface7fcad1c494c2ee5e7176a2e03;
        49 : storage = 256'h02788a5d58f72cc9210c30d50731827108d184a5d56e655bb235156305717e67;
        50 : storage = 256'h4f8038d92e830053b8869cb7afae17b15aed7dfd37e0a65fad5381969748b483;
        51 : storage = 256'h24c75b34ec81340644875e60823f88215925bd6c2e2fd691258362acf70d21c3;
        52 : storage = 256'h19e3756ecac381d08571c906102864c123b1ec524bf96eb171a7d224ef7e0bdf;
        53 : storage = 256'h1e27ac0e70e98c9a590453a7eda612e151bdd845da3db481bccdba0ace4adccd;
        54 : storage = 256'h53b5818e11a2dc3cef7f24d5a05c9c01554e5e94867d00856de7157a82fc4499;
        55 : storage = 256'h3a81de5228ebe73426698f45ebf5a42173284539f4f5c09b7f82dcdbfaa4dd05;
        56 : storage = 256'h048c4be581c9a51af49aee928dbbe7d15d7767f10b171c63ef81412c5f8ad17f;
        57 : storage = 256'h008ad0c371d6b9a3b871763fe0162ea10207d48f36df01bfd4d86370331e92e5;
        58 : storage = 256'h263123f9db8443e287a1fcaeb69ede914e5193eefb6d57e42ba2d61cd89450a3;
        59 : storage = 256'h467569a4d1f30fe3e15493e1ad3f124160c7980d3d5a562dafd1cb1ce7444571;
        60 : storage = 256'h0f725f380e13cd608735ea965ce368f173ebacefb5c5c427dcdc3583b964fe0b;
        61 : storage = 256'h07a91bfe07a3cab5a6c253948c32700112c4527107ac4573aab12a04f6c894cd;
        62 : storage = 256'h121af97e39cda196ac4078f6e703ae79135427dad0f2a61df4fccc56b486d923;
        63 : storage = 256'h0fc47525f3531fbdb333f1637bf44f0110c0ddf9ecfa913d185253c298146b0f;
        64 : storage = 256'h00b7be3991cf9158ad55bd25c9e587d1017f9fd76b30397b7cbf425b89bfd043;
        65 : storage = 256'h0259fba90a47843f478aa01f1ca7620d0edcd18931f5a4c581b179ddf6f0bad5;
        66 : storage = 256'h1552ca2fc02327e15fc7e792e4979a791f0b966a7fb4281ce64a873f7f345059;
        67 : storage = 256'h075d01e90a21ccc0ddf611da7a5dd2490af0ac91119ff4512dcb206ba1e52b8d;
        68 : storage = 256'h003443c040c8a69c4a38ebd5370a9a09026d31e30de096487adacf27e1d4d199;
        69 : storage = 256'h001591e0822b742d93256bd20f991bc104322e5027ad32c752821d9aa807cbff;
        70 : storage = 256'h0b1f7d3727f9ad90c45f20ae10ccd7a91ab982cebac1249e9e595e6c70fea83b;
        71 : storage = 256'h0104a2ee5e24f216294d153316c3349103c8ef0287209aabd988ab262340006f;
        72 : storage = 256'h10319ac2a8b5b89111ea1b3e02f2d0691719c5787ae74cbfa8e6a5afe6d988dd;
        73 : storage = 256'h0d67d4fc9bd3044e63e9698239a1039d17079e7c4c4185c2a51b7602f702e705;
        74 : storage = 256'h01ee62275c4c59d0ece4a1a274eab67102c5d1b4ff0005e8726d78b245cc279b;
        75 : storage = 256'h01f42d0faf9e2f6b872d01d44a49ee8507b28bd312e9511d1b8433f0da33f675;
        76 : storage = 256'h03198ab43d875dbdc9ef49f87e8ebcd9053252e704e0448ee9630f4957b76ef3;
        77 : storage = 256'h13822f0e1b7a0515476382890c7b316116da8fcc36121641fd9f1280fa7fba45;
        78 : storage = 256'h0c54c2d164822eb9b509a4dd69269f0113a7f9c30cc969b79dff033d09ea57e7;
        79 : storage = 256'h01362eb3f437c1d2c917549958ed57c112ba70ac218d68015f9a0c7c13fe46fd;
        80 : storage = 256'h02027dc99598ab4c4d7f01cc662a8711021154130bfc35b65fce9748087e3299;
        81 : storage = 256'h003a368e0b8bc04b5b03ea4700f8aaf51551f51b81350bc303f51594579d407d;
        82 : storage = 256'h109cd24ff2aa5fbb74e5bb03da809ae914e718786bc95178efdbafe6e6fd933d;
        83 : storage = 256'h02397ac293ca75659b5cb256ba178aad085e9a0cf0ebfc6aa03e25f221eeed21;
        84 : storage = 256'h0355c88042076eae15e4b32d002d47a1132a8ee815012ee8ad3588efea925e33;
        85 : storage = 256'h12c9b688e505831623f07ee36265d5811400856b4b64a6bec63156990dc90a67;
        86 : storage = 256'h0a9bcf1d4508a3cf2177dca06ba4d9691b0058605c525e78c04045724bb0e5fb;
        87 : storage = 256'h00fe13f22d345005592d9026ff3e9c6115ea58586c3433e601df5276a33d8781;
        88 : storage = 256'h00398b60363fb3e94625f29baf863de90079e2f0bb5181b35bc0b50805ac501b;
        89 : storage = 256'h10f46db36841849806ab45932e39076d125d18c53f3dc6f3fa576272175a845d;
        90 : storage = 256'h148c89fbbd158c3983d5752a5310343116b139080ee0febe751fbce54e51f18f;
        91 : storage = 256'h193b94c4dd5ee5737decc68858f9c72d1b2e299dace15bdf3742ba1bf8c4aef5;
        92 : storage = 256'h015bc6b1949d69c5ee5a4905b38538b904667c983a307065fdb94ca3591ca633;
        93 : storage = 256'h06a80e748815568de2f7f64ad6016fc1075f9cfc07ba357f68964987448cf1b9;
        94 : storage = 256'h00c2d3001a2af8d6bd12674d4da1928106641be9dcef6f327ff5ff80db8cfabd;
        95 : storage = 256'h00b7be3991cf9158ad55bd25c9e587d1017f9fd76b30397b7cbf425b89bfd043;
        96 : storage = 256'h0547d65ecabe834de09faf0c685beff905ab74801fcbd9fd26ea454d62471eaf;
        97 : storage = 256'h07d51b321bdec0076f1092db7bc278890bd7d4b6a4a9b999e23f08e375fe7cfb;
        98 : storage = 256'h038a7b91b346dacb4a38a3f973e9dfc9042c655c40960aa0c4ee200853901957;
        99 : storage = 256'h00dd547fdf695907fb798f50af08672900ecf8e63dba10f1b5ac25faf6c0ccbb;
        100 : storage = 256'h006657aff9b8983a088d1bd9f8b9a6010199c6caf8605fe2a9b40133cadfb68d;
        101 : storage = 256'h08769daa79a7f72c85827a46fd6cd7210a31e309f67810e37c14b22f68b83181;
        102 : storage = 256'h003c5a7629088739b06c71dffe7da4610171a082fd812a9cda95b2a913eaf4dd;
        103 : storage = 256'h086cbbb55406767f46cc9371ce0da93108cff9788ef52ebeba532c683a791447;
        104 : storage = 256'h009608f7ac043eef37784dbbbfda67a108c90cbf69dc925b8e79229d2499683f;
        105 : storage = 256'h00b8660d19ae53911bbac1d2d0aacd21010ec7ce87df4fc9280567c6f27449a1;
        106 : storage = 256'h00dcd8b9ac6da812c32fd7d022b07fb102efb8651e1ea3f8e33a5d7a992e078f;
        107 : storage = 256'h00b1381299ba2bbef467e586497081e101fb7d4d5bfa9a3e8a606bc09ed1ce29;
        108 : storage = 256'h088897d3de8f3417e8a880509a1eaf6908b7dc8436b787004bc8f07f983e8dff;
        109 : storage = 256'h0690d0bcaf67be15702d3e8693be6101077f96b4fcbff0dba5477287038a57c5;
        110 : storage = 256'h058db125b3a11306a626e263922bb2190724f95e61f4a04e45fed7be9d7e1ca7;
        111 : storage = 256'h00a85af8cf4e28d64bd6435ea053907900c9ed5e36ea0a9e7b75a2fa1fa45fbb;
        112 : storage = 256'h034dc5f0d21676ef6f3319ea05602031082217694bf0ee89fb2e691404e3b127;
        113 : storage = 256'h024824cb642ec3294b81e722d5d93bd107f95373cbd4873283242b48aec49d67;
        114 : storage = 256'h023a6dde0783ee7e53be6aea1fd0df7103315b113c50686eec1de0f503d812d3;
        115 : storage = 256'h0099da76da64deb17294c0c192db4d71074fbea4c05ae9d32fb1a94b29a987e9;
        116 : storage = 256'h06db3091f553c6e133b4ca63261bf80107a15dec33c64092717fa81c61d50745;
        117 : storage = 256'h051024cd2c12be80c9b3e8ee02f7dc210a4ce89959770c69abf46b3f92f4aec1;
        118 : storage = 256'h020a79996955f1f96c756c0aa673a0a9085c39588438d313f6646158a5924bf3;
        119 : storage = 256'h00021ae2950db86e2282d19a2bc316d1002e7f3d576e235d11d5c81e47a4fb21;
        120 : storage = 256'h04011dd696055b93d7a12db7fa884af107015d9ac0a6f81feb3468493f3f8ec7;
        121 : storage = 256'h02dae5b6bf8f062a241bdb124d46aca108a8176c28c35874012b5ac8d4b4e63d;
        122 : storage = 256'h00b7e12caa62cccdbb071d9edd3df1e10a5e630c27aab237ede1665aacff690f;
        123 : storage = 256'h019165a14783c99fa18cd0fd56057a0101adbae47ce05b25b3e336f6b66fdfe9;
        124 : storage = 256'h17dce7f8240f812aa23455c8273892094921813d53ecab68210ac49ed1d7870f;
        125 : storage = 256'h2c2800c5b77cc50180cf51483bc2e3213f6310c0d9d99a749bf589b203c9d22b;
        126 : storage = 256'h0259fba90a47843f478aa01f1ca7620d0edcd18931f5a4c581b179ddf6f0bad5;
        127 : storage = 256'h0547d65ecabe834de09faf0c685beff905ab74801fcbd9fd26ea454d62471eaf;
        128 : storage = 256'h3c32106d05af53604dfcab4ec0a3dab97575f3764c3992365b35b83bbfcf9bdd;
        129 : storage = 256'h173ced3a6437e11cbbcfe34f724832f529647092bcb2da8da92a52d3e1b0f661;
        130 : storage = 256'h02853c3f30f6251e29c998cd184b10e1092e4f83e329dc8c89dc23ea069f0a1d;
        131 : storage = 256'h0b956ffa0f2a8565087e8b5e36f88ff10fe0329ec526dffb05a40d9fe32c64db;
        132 : storage = 256'h2528d3454675922e0d96df073b1f3cf9651d132fbb68c6ef148792c669839d87;
        133 : storage = 256'h0c5c826f60c826b5df9fcfde38f190410e51fdc5e930da1276d034726e82090b;
        134 : storage = 256'h07243f35544c13ef9c7373aa8a5d29fd5766f14da928064cd82a6fb8dbe4a2f1;
        135 : storage = 256'h22b8325b9c5321bc579c89d1e97c9a49572243497dc329819221ccd14c94d6b9;
        136 : storage = 256'h014dc59551fb9b9b3b6ec0938be815d90a7d9f9b286ac98f505a59fcd4a8a667;
        137 : storage = 256'h0a04c4065adecaca84179fcc88f275851d1f9fd5d662a6246bf976b4d28f21e9;
        138 : storage = 256'h00e9efc2e9b343a0bcd8090feab381f113a9529a6dc6f615d9f8a5d337d2de1f;
        139 : storage = 256'h527dc71a041c8b0216f63ea699a72fcd5677c96d81061c07aaae244cae9a1ef9;
        140 : storage = 256'h29a31afa9fa49aadbac9fb835e693a014a5ea3ea6ae1d9015270263b64bc7563;
        141 : storage = 256'h3e1ee8abf60993a1a7bf5d86fe378a0d46dbeac93886e3a3f374e17c4848fd91;
        142 : storage = 256'h06fb98dc5fdbeeb4494dc1496fa4373d07d2bb1f1446d64f62ce52851cd10f1d;
        143 : storage = 256'h46ebc08246be0d96e005a6087c9c761150aa5b28da8569b6cf3cb0b502ad8d11;
        144 : storage = 256'h1a5a00bf758a3db9bb100c48ed4b23a54f160a7368224525cbab77b96908c2d1;
        145 : storage = 256'h067788d2e8201fb1cb48be000877e0611faa9a22e808b7f7c2f0c4c2a91e3cc5;
        146 : storage = 256'h414afcc7772e3d57bbef64239788daa948841e9abf6c3d334fe1a6c0a6f6325f;
        147 : storage = 256'h15d237c73f4570cd3db7f47855742f814bada7b83dd6a0ca719ee7e1a9f5c1e3;
        148 : storage = 256'h23252aa90a35876eac55ab11cded38b16629141f64d5c1c8d133429626d2ca47;
        149 : storage = 256'h096cff1a2b89abb8c408ff9c64d19df952eaeb6c31e385c20fe02a9a34592ca5;
        150 : storage = 256'h00bc33d2c5d0ae2121e9b4b378fdfbf101cd2951edc544c30dd668ce97b200e7;
        151 : storage = 256'h450581327e2528df24e36a9b16ac4435457abfe10b398ce9957bcd4bb1217c71;
        152 : storage = 256'h0c9f531bbf2dccff1052c2d9d74c551155db6131b83fe0e3467107f635c3c2ab;
        153 : storage = 256'h26e1ce6e9f75b40238eb5fc45a38fded66d66e130cc3371f3e9c7297a20d4c69;
        154 : storage = 256'h073c7a73010f35cb630d6a6b70b1234910a6192d6d01ec052e38018a4d6a9a5f;
        155 : storage = 256'h381a8dbcda8291a3355870504867ac5198c1e2da1e53a3eba02ec1fe860b90db;
        156 : storage = 256'h061546a164f2d426653034353f2806f184677269388eee00173730535af320a7;
        157 : storage = 256'h1552ca2fc02327e15fc7e792e4979a791f0b966a7fb4281ce64a873f7f345059;
        158 : storage = 256'h07d51b321bdec0076f1092db7bc278890bd7d4b6a4a9b999e23f08e375fe7cfb;
        159 : storage = 256'h3c32106d05af53604dfcab4ec0a3dab97575f3764c3992365b35b83bbfcf9bdd;
        160 : storage = 256'h3c5afe39c781ab381303f932b676dd9d567612d6f14645199dcf26027c8bb355;
        161 : storage = 256'h06ccd5a9e8116ec4831894553b86c69d132d613eff521c78011fa9d369e19441;
        162 : storage = 256'h087299706560e4ced01084ff18ebc751212962719b36e9e755400b2fac515b17;
        163 : storage = 256'hc9d5533c35900b8811312d7fad68eaa1d3354e9a6ae264cac9f265eb45768db3;
        164 : storage = 256'h1c172945fcf29f2d191a0e582021b5911de99a2fe7030cab423a03fea9ec1507;
        165 : storage = 256'h85eba5808fede7706e31a61acb5a5ff9b691442c6065db0a9bee1532b14da125;
        166 : storage = 256'h9a3a21aa91a68b132aadcbd7dd75a809b601ce79c4deea100f17ee78eb78d38d;
        167 : storage = 256'h048fb7d0fc9499327f96dd3b8a7f099115e9c9e4af4cdc11e527eeec97ed7c13;
        168 : storage = 256'h00c4c1ac8b5e2f04171eab9c4d6027113cd5785d1364e935d2f76f73cc02e07d;
        169 : storage = 256'h0c9886363201a143c4306bf30986c1612911b6b9718e06b2323a288a1cc4eb2b;
        170 : storage = 256'h35b31251dea063a0723f6b10c51000adb49db6695afc781a0e73035800d918cd;
        171 : storage = 256'h9340af888fbef1d7e214b3c0345d66819b58535868f6e53633857bdac693313f;
        172 : storage = 256'h01cfafc0e56d7f2ff528063fa96ba29994030d97adc576933c41f8c04608ac45;
        173 : storage = 256'h01ecd88065d699f9db5d4e0b41cdf72510575910e3495e6a53aa4903af5add41;
        174 : storage = 256'ha382b5556febc510037b490ee38a4a29a87ee99ca93a507264c59d061231c1c5;
        175 : storage = 256'h7fd91bb6b0d0c1a04d659dbd0632a981a5325eba20a9d832d074a0e4cdf91285;
        176 : storage = 256'h18f28f634dcf58491efca8d866b3271942253f2240879cff9958300b9ef72309;
        177 : storage = 256'h767293878e17864a152c577cc1357881977922e5df62cf2e1437e269db8cac6b;
        178 : storage = 256'h1894ca0b711119f83dbb2e8f5b6807819e141ca490b4bda5b6675c0f058ba7bf;
        179 : storage = 256'h000e2ba8d9d1f8ec08d20a5ddd13f869d5651e70a2fc1e3a3013dcf8153cc173;
        180 : storage = 256'h8c0b37b50a8eaa47743b2a0482fad72dad33403fb3f5603776038d77885fa469;
        181 : storage = 256'h001996fbcbed67637ad43f64826da80903c348b20dff9af80e73ac36a31a5893;
        182 : storage = 256'h3232119e1161c3a6e883cfa10a4c9e45912159534ddeb1cd95cf04e2c5ca88a5;
        183 : storage = 256'h8a1186e76ed9e89dc4721761db692c31b35701806c23e654d6f70017607a8b27;
        184 : storage = 256'h4ef598acae1c11c3bf4b4eb021f29f99d6cf3811ecd6520071d1e40422e2ccfd;
        185 : storage = 256'h11a187b77d182b694f344dcdb0a0e07122c6c37e88dd981fc5b07de0a5e8346b;
        186 : storage = 256'h03008bee2c7fce6a0872306035c1c25935d4a3ce70e79ea2ab62c906f429f2b7;
        187 : storage = 256'h1c9df7496f3019daeb9734af5408edc12ea884849d310bde5d17b981f6015973;
        188 : storage = 256'h075d01e90a21ccc0ddf611da7a5dd2490af0ac91119ff4512dcb206ba1e52b8d;
        189 : storage = 256'h038a7b91b346dacb4a38a3f973e9dfc9042c655c40960aa0c4ee200853901957;
        190 : storage = 256'h173ced3a6437e11cbbcfe34f724832f529647092bcb2da8da92a52d3e1b0f661;
        191 : storage = 256'h3c5afe39c781ab381303f932b676dd9d567612d6f14645199dcf26027c8bb355;
        192 : storage = 256'h0418bb17797a22f8232272e150bd6c4106c207f0aad9506f65c9bc1da2246795;
        193 : storage = 256'h0838f154d15189fdc5295c2a64f5fb110baf997bb2c78da2af28a5561762e0a3;
        194 : storage = 256'h4121235b574ae4e50b9b3b9d9b1681594a6da4f726a767e915bd9a61257ab66f;
        195 : storage = 256'h05684311875b462d093b1705381d9e110a8a7c3d937730a3b84a6e330a83bd53;
        196 : storage = 256'h14e7934adb43a1771a74eec48ecb01fd4055e27aea6105ea66576fc9e06fa749;
        197 : storage = 256'h1ac5a49edf23422595c88fcac0b21eb14023549a1b5876f8df7477a2c69a13d1;
        198 : storage = 256'h05f534d603e3d9a902360d97a90ed2e107b8d9a3bcd094256e6ebbc726bd1c4f;
        199 : storage = 256'h030654df9a1b6b7686c3d8026568a02d156ffb4ab15220e3e2926b27cb9b7f81;
        200 : storage = 256'h0c06a3283717e2ea451e9534ca6ee3510e78f57e2c2b7bac583a24022d374f47;
        201 : storage = 256'h25af78db5925d4ae5cbcfb764c658e113fa5d86f5ffc14827ca18977ef229211;
        202 : storage = 256'h33da6cc9f2abc119d5198fef7609730136be14311efa228d37b48540b1de2beb;
        203 : storage = 256'h18636c85f967eae4bb26dbeb244734d134288a8def12ea7d3a0db0d8415a18e9;
        204 : storage = 256'h055ba1fdd0a2e617727febf219ca849905c22eb50e44c302d6d9532e6d07a495;
        205 : storage = 256'h24ac919a87bb9e0a3d6d79b8ed7253fd3b6070c4c4e017b8151e0277f69b3c69;
        206 : storage = 256'h17a668d8e2c70b8a122436fe291295053a36d4639ba82def9dfababaa42b8c29;
        207 : storage = 256'h1008ff9d43819c8573521c8f5211656d174f2843edb5bdbb9e4afebc58a8bffd;
        208 : storage = 256'h25517d555f9884c6cd35083c1e37f9993560ca6ddc5a6173aeb6ebc30363f987;
        209 : storage = 256'h32ec421e6c17da11ce515fb9fcd4c10137b4adbcd6318231c6a2e2fa33e8846b;
        210 : storage = 256'h3840f4f92a0fcf9fcb247ab930996ff14b32eb0d14a18193085a519162f6652f;
        211 : storage = 256'h38990b2fbdd0bd6a70564cfe0c059a8d3d08d7460d5af6a73d471c28380af4dd;
        212 : storage = 256'h0007a5233665d7f90b26ed54e5134ce10153745acd89c6eb652ca9f4af8152cf;
        213 : storage = 256'h2858e86ab23fd2dca4c08bedf289b61d33249457376c5102973c8b77a64184c9;
        214 : storage = 256'h09ebfb701cd9775c7ebbcd5622b8cb713f32b75ff9129760fa9d1207d75ab5f3;
        215 : storage = 256'h08808fa303fa0f1db36e828ed5c5dc554bb2850ba31c61cab07e1dfdcbb40601;
        216 : storage = 256'h06a93bc1f8966d9ead0d5f6050b338b10c41457d08d0485d3d0b40213a382187;
        217 : storage = 256'h04a4eb17d043e79c33d1516294d3be610bf0928161207ef073aacfdbff82789b;
        218 : storage = 256'h056b6af8b956690804a7d01c1f1945510a59511e196dbf33ac97eba82ce1df67;
        219 : storage = 256'h003443c040c8a69c4a38ebd5370a9a09026d31e30de096487adacf27e1d4d199;
        220 : storage = 256'h00dd547fdf695907fb798f50af08672900ecf8e63dba10f1b5ac25faf6c0ccbb;
        221 : storage = 256'h02853c3f30f6251e29c998cd184b10e1092e4f83e329dc8c89dc23ea069f0a1d;
        222 : storage = 256'h06ccd5a9e8116ec4831894553b86c69d132d613eff521c78011fa9d369e19441;
        223 : storage = 256'h0418bb17797a22f8232272e150bd6c4106c207f0aad9506f65c9bc1da2246795;
        224 : storage = 256'h0000a8799ac2460a5b9a604293d0553102978ae169dbc378e5a512bb1ec805d7;
        225 : storage = 256'h0b371e11c474c76507f4ade725be0be110822280da9e589b01f899a581e43373;
        226 : storage = 256'h00cf9d0ccf3c012611ae25a72e3869d102568779fed0c3849485fb5cac590bc7;
        227 : storage = 256'h0282cc10164e2d516c445d67ef97e9910e450d4b70d259adba0bed7480793965;
        228 : storage = 256'h0a6e0b6fd0ee65cb3b48731ddddc6ddd0e39d6c2e830d6e0095ecd8409ff3dcd;
        229 : storage = 256'h0079094049ca53307b452d0f8161aab901b67819f7932ab464bfe21c6005d9d3;
        230 : storage = 256'h03ec0a706df78f5cd5b566e2b8a2e05904c13eac83289c1bf62ba243016d56bd;
        231 : storage = 256'h01efaa713b6b315ce2cfada561e814710335c45918e247a0865c44cf299f56eb;
        232 : storage = 256'h0132298fa9c1c9a8f74abd9812868f410e1e018f46e41f7c0bb2fffe26b8930d;
        233 : storage = 256'h060a8ffa168d3631a3fd0390a470d0010c245979247c34c0562edacaf4e0ddff;
        234 : storage = 256'h0a4e036bc687a2efa5f9ab441ef880610b919e832efdb0e333925cc0e8846c85;
        235 : storage = 256'h00d972e5caae9aa3f162c860c4ffe9010146f9fb194e68fd94b840f21d2c5081;
        236 : storage = 256'h04f0cd7d414c5afd0af1cb7226d8f2790d2b7c9dd6fde651d1be84caf9436205;
        237 : storage = 256'h0b0b62c147582ea9bda2a06724cbbcb90ce979e362b16a922d6089bb229922c5;
        238 : storage = 256'h0113d8521bc446b944b47c715e9d0e9d052b86e30b7f067577f79588d4a66049;
        239 : storage = 256'h07f259c209c8efc11bc346323d2555b90bd6e0713f5a381aae2410462693282b;
        240 : storage = 256'h05039dcabbcc4cfb202a14578663b2010c5b0bba2c30e7b3d469a28f28ca747f;
        241 : storage = 256'h0090820892e7d7eb19287018977e0e1110ade3f669c5b165778d53462eba9733;
        242 : storage = 256'h00517d1653239a92ef6a72bc88b17aa50d899e9e858da860c9634f7c2ff759a9;
        243 : storage = 256'h003da83e6f6d186888ffa0123dd33ec9004b4aaa384b057d24ab8067acaf5653;
        244 : storage = 256'h0818143a9f60673661b0aec2b6ea6e450b57f58c36c85849893320078cb680e5;
        245 : storage = 256'h098ad57ff2f49b0340b656fd1f2d33e10e047860e86587a9a3df0e989b7369e7;
        246 : storage = 256'h0c232ef27923f1b23cfac2c95ca9c93d10ca3157b441a819de6e5b9c65bde33d;
        247 : storage = 256'h00b7843866d9f79abd9959ec27aeff6102b7da51913ef4848745b63c3d68b02b;
        248 : storage = 256'h117e43a455df08211532593ff4ca610114a57a46db9cd9e76da1f1aa2d45ffad;
        249 : storage = 256'h023e412d8bbc948e1ca4df15db1f924111e53e99690d80a1beeec0c112f75b01;
        250 : storage = 256'h001591e0822b742d93256bd20f991bc104322e5027ad32c752821d9aa807cbff;
        251 : storage = 256'h006657aff9b8983a088d1bd9f8b9a6010199c6caf8605fe2a9b40133cadfb68d;
        252 : storage = 256'h0b956ffa0f2a8565087e8b5e36f88ff10fe0329ec526dffb05a40d9fe32c64db;
        253 : storage = 256'h087299706560e4ced01084ff18ebc751212962719b36e9e755400b2fac515b17;
        254 : storage = 256'h0838f154d15189fdc5295c2a64f5fb110baf997bb2c78da2af28a5561762e0a3;
        255 : storage = 256'h0000a8799ac2460a5b9a604293d0553102978ae169dbc378e5a512bb1ec805d7;
        256 : storage = 256'h0c101ad9fb7cc61fbc1c53649ddd34411c8be7c36b32f2dd1c68d3c3e0ba9715;
        257 : storage = 256'h019d08de44010891b6f376be355f5f81040afcaf4b93d3a0f303d8451968cfa1;
        258 : storage = 256'h0b4b08c83bc595f96262bc8ea3d7bfa118aceba9cd0297ade73beec32ee57e53;
        259 : storage = 256'h10ebcae521abf6f5a3ca08b9f15d3781189987e32d7b64757e6d01c44ca825ab;
        260 : storage = 256'h013d89f5322b7d74d76a0869a372252102f6355b90a42723ec2cc968274581b5;
        261 : storage = 256'h014384dca78c888a239b60f7318898510838e17b4bca6db519e1d9853bc80f3b;
        262 : storage = 256'h01ce45fd539233703f24c997c6ce7901058d03805addfb9c9deb7a73754d5cdd;
        263 : storage = 256'h086d5a756222e70d85bb7cb787ca9e01186966dd90069f25ee621cfab87f5e6b;
        264 : storage = 256'h11946794d964ca7c655f829a55eb7a0114ff02ff0eb7a78447e374819793b8a9;
        265 : storage = 256'h0306caab340c31a33a6f14f6a517763114014879a0d05adf5715daa34a45fe33;
        266 : storage = 256'h0112510a036a66523f80c142b729fdc1023569d44d1214c745f1e7b61a0194d7;
        267 : storage = 256'h082b0b4e34504fe463075eb9a1bd8c2116c6088229c2d6dd7c1b12ffa614ecb3;
        268 : storage = 256'h071bf09ef11f3c0f7099e1abcdade0b11653e2ef6c2bb070a2e21bd2de442df3;
        269 : storage = 256'h03fc57db338a43e2f17e854f85eaade108f0aa64dc127feeeb817dbde2cc79cf;
        270 : storage = 256'h045f07efcf54e75222db201f2ace252114790b6061da9e042debc30bc4a0b99d;
        271 : storage = 256'h0f4256ff08661480f7f93282587f4401155d97efa1ddf6a7f42d2f5e1a385e29;
        272 : storage = 256'h1aab3d9492b73e4784371e6d7273dc211cd7918531fcd5fa42aef38cae6c3d55;
        273 : storage = 256'h0e2f0e2310cc69ae63a6ce006194e3311768cf30f8620247171f82fe4667996f;
        274 : storage = 256'h00792b257f9921e7ad342063d6d777e100823215758fe6263207e1b3be575135;
        275 : storage = 256'h129837ff861d2d66bf007c904a3b21e1139d938f48b314f192e2499565e44ad3;
        276 : storage = 256'h03649f5ed0e5b7cc03444799da8ea281183d3ea8aa3c2eb56c2f85b9a803ec81;
        277 : storage = 256'h0d7c85693c89ba430c9c1cafbd4022f11d08825b52b2030558239329e7304ebb;
        278 : storage = 256'h02e93ee28fc7271258cf13225dd2b1c104b347dc44d51e32186c85f37e79f19d;
        279 : storage = 256'h61712f61799db8153872bd75f36983c1837f7776bcf6f6988de70714dcc3d721;
        280 : storage = 256'h50bb68596a762eb1136709a1dd3386a171fa2bde6b6fa15e4477bbcbd1ff5ac5;
        281 : storage = 256'h0b1f7d3727f9ad90c45f20ae10ccd7a91ab982cebac1249e9e595e6c70fea83b;
        282 : storage = 256'h08769daa79a7f72c85827a46fd6cd7210a31e309f67810e37c14b22f68b83181;
        283 : storage = 256'h2528d3454675922e0d96df073b1f3cf9651d132fbb68c6ef148792c669839d87;
        284 : storage = 256'hc9d5533c35900b8811312d7fad68eaa1d3354e9a6ae264cac9f265eb45768db3;
        285 : storage = 256'h4121235b574ae4e50b9b3b9d9b1681594a6da4f726a767e915bd9a61257ab66f;
        286 : storage = 256'h0b371e11c474c76507f4ade725be0be110822280da9e589b01f899a581e43373;
        287 : storage = 256'h0c101ad9fb7cc61fbc1c53649ddd34411c8be7c36b32f2dd1c68d3c3e0ba9715;
        288 : storage = 256'h15e794f0ad45ae891dbb4b5d2bc5056119bfe222c53b0957b791998d6b3df9e5;
        289 : storage = 256'h76ac64137c7356c9907fe30a773d41819d28c6f8f7ad003d0936a07e608e1edf;
        290 : storage = 256'h56fc96358cf85dd41ff23f1b6dd708b19cad4870b4a9537eb096286793526d97;
        291 : storage = 256'h10c05e85391d1dcb0572fbbbdbc3af7112dd11140f94e9c95186e790e0b37f49;
        292 : storage = 256'h1e0fdd5c1c59ff328605373eb15c6c11345e16cf01638c15f85585f1b16ad967;
        293 : storage = 256'h1d7c243ac2b170d82fa472a8b73cd5e1235a8181f77ed27ee31ec51e25951d11;
        294 : storage = 256'h889c0653bf0caf00a68ecc6494401aa99b7abf3f1d172ac698eea2c28b175957;
        295 : storage = 256'h10d2d574d87e7927459fa642edd1770185b9b6a6eb2517c018e5ffa519f8e50d;
        296 : storage = 256'h01e83e26f87e35196b78b80f2ceaca997f69b41deae8ab18cebcfb8a36a6263f;
        297 : storage = 256'h0318d94a31b6b6a869016318204198c90e11254b675d104afe2569ae298c3e73;
        298 : storage = 256'h1b7c52660614aec9d3d5ab750f0422a9910bc4994adcca1219e908796cb72ebf;
        299 : storage = 256'h72c27173ed83bd6bae9162cdd15889418e34c2f6d14c4c990bae2367697c24ff;
        300 : storage = 256'h036853056fef90edb917f58749d8529138f09fa449f44ead4c3d98e98dc2d94b;
        301 : storage = 256'h5125d9aaeb4ac833548a8830c964bae18264782a4f8c6e4ffc434cff9f8dbcd1;
        302 : storage = 256'h2d654002a5c727f78aee0213bd86bb0188141c0de27d8540fbc129ccefd4c08d;
        303 : storage = 256'h11b1ea74d497f0df0d16493d28825411b7b24f5936fa6c3cd0f473e38e76c169;
        304 : storage = 256'h87bf94268e79a72d7eab95dd687475b195187f395adc2ef4793ea27911830f6b;
        305 : storage = 256'h020a3429ae4e487604348cdb17da1381033d38f0c806b0fb6da37e59e52eacc9;
        306 : storage = 256'h2f66d6f78549fb221524d71e5ba1fe717ceeaaad5f9dd45ac96f765add6efd5f;
        307 : storage = 256'h0ad393c1e8bc28ef29838fdeec0096819a6182330c979941a3948b0a9f57d245;
        308 : storage = 256'h3c15963760c9e57d185537697f985ae9b8ea041f7c10f42d625b2a5d92ba36e7;
        309 : storage = 256'h19a829d8a72a394b9112d99f647c09811defc0ff4fd41a106a6e0ff828ddd4d1;
        310 : storage = 256'h0b379c19021b0a33f958243fd67933c1129f9c7e6ce6b24a30f2a165d54ebffd;
        311 : storage = 256'h039da2740844df6aa3a8a4b4140f0e01102460d94389d477903bd88193721691;
        312 : storage = 256'h0104a2ee5e24f216294d153316c3349103c8ef0287209aabd988ab262340006f;
        313 : storage = 256'h003c5a7629088739b06c71dffe7da4610171a082fd812a9cda95b2a913eaf4dd;
        314 : storage = 256'h0c5c826f60c826b5df9fcfde38f190410e51fdc5e930da1276d034726e82090b;
        315 : storage = 256'h1c172945fcf29f2d191a0e582021b5911de99a2fe7030cab423a03fea9ec1507;
        316 : storage = 256'h05684311875b462d093b1705381d9e110a8a7c3d937730a3b84a6e330a83bd53;
        317 : storage = 256'h00cf9d0ccf3c012611ae25a72e3869d102568779fed0c3849485fb5cac590bc7;
        318 : storage = 256'h019d08de44010891b6f376be355f5f81040afcaf4b93d3a0f303d8451968cfa1;
        319 : storage = 256'h15e794f0ad45ae891dbb4b5d2bc5056119bfe222c53b0957b791998d6b3df9e5;
        320 : storage = 256'h0b55ba6c708dcd5c500e45fc4b7093d11641fe8f2b06733e951daa2e20bd9e03;
        321 : storage = 256'h0265d76e68e11a152aa1c2d57f0d7c611630812131f058b85bca878560ab2edb;
        322 : storage = 256'h01f503baf4c64d09296e422133586a4102abeb7b406e3cc3923cfe186e11be85;
        323 : storage = 256'h055e4eb8a2292817324478e463dc8121076aa57ea3b2637e571f857f096fa96b;
        324 : storage = 256'h03e070bef1c25eb620c72ac3e9d7cda10501c8b6a48b969a535bcbe483b3982d;
        325 : storage = 256'h117f422294915e573434e6ee19c533411605174f7440323a12d336ce13e2939b;
        326 : storage = 256'h00915e7b6031698a61cf6f8b5ed2d60112f05f764075ffb72d4034f3890d5ab9;
        327 : storage = 256'h081e4ee8e73e740c1d839bf53249f371120b81204ef82756c1d81cd46a14abe3;
        328 : storage = 256'h01b0daf4cf474c802ea4b7bd34966a6101fe03c3679592255e6865442a980ac7;
        329 : storage = 256'h0173708c85785f2d20d86de58aca72f1148acfd4170e3faf62d6703d80c94263;
        330 : storage = 256'h07ce655f5c46b2db194dc9f21cdb84e11423d95bd3a3318b4fc2e8f7a57af7a3;
        331 : storage = 256'h037703223b40eda26369ab29d4274cb108106c98d3bece467c7777788e66633f;
        332 : storage = 256'h118e1a0dad63fe32cdf6b99235b977e1127788189622e69fd1e4fcbcefc760ed;
        333 : storage = 256'h10d1b1a7b94c97743650c1fd91ccf6011345b00a258de98bdfbbb96ccb2b9839;
        334 : storage = 256'h11aafae2c8bfcf78f2e8b8444e5ac7e11a04220fb93e55ad513bd5e4f1a1e425;
        335 : storage = 256'h113536496217892dd991a58963ecf201151da3a7c45668f1cab703251a2f2cdf;
        336 : storage = 256'h00630756d6deaca31cbd209d158e35610075706ea67c6a20b01d0ac893d2c605;
        337 : storage = 256'h05aaa5bc696e39c6382310117e86917111b1911e7844d454c854ab83bf18f283;
        338 : storage = 256'h0216d0263c44c68f27cf3ec02573638115dd42ae023fba2cc1ba670d17910011;
        339 : storage = 256'h154ad3749fdc9aefc59ecfc8a94ca1c11a304755705f4b91e6800b4ac2f620eb;
        340 : storage = 256'h004c3b6be863065de6ce757f16d1e121043d62646e814b141127cb78353818ed;
        341 : storage = 256'h27deb6f076fa39e40de1ca00741e69e171aa8ca9f5dfab875f0cfc77d4d373a7;
        342 : storage = 256'h26b05441fa797fb114f9814623e0f78162857af844b5b2489ab99e11d9e5cc23;
        343 : storage = 256'h10319ac2a8b5b89111ea1b3e02f2d0691719c5787ae74cbfa8e6a5afe6d988dd;
        344 : storage = 256'h086cbbb55406767f46cc9371ce0da93108cff9788ef52ebeba532c683a791447;
        345 : storage = 256'h07243f35544c13ef9c7373aa8a5d29fd5766f14da928064cd82a6fb8dbe4a2f1;
        346 : storage = 256'h85eba5808fede7706e31a61acb5a5ff9b691442c6065db0a9bee1532b14da125;
        347 : storage = 256'h14e7934adb43a1771a74eec48ecb01fd4055e27aea6105ea66576fc9e06fa749;
        348 : storage = 256'h0282cc10164e2d516c445d67ef97e9910e450d4b70d259adba0bed7480793965;
        349 : storage = 256'h0b4b08c83bc595f96262bc8ea3d7bfa118aceba9cd0297ade73beec32ee57e53;
        350 : storage = 256'h76ac64137c7356c9907fe30a773d41819d28c6f8f7ad003d0936a07e608e1edf;
        351 : storage = 256'h0b55ba6c708dcd5c500e45fc4b7093d11641fe8f2b06733e951daa2e20bd9e03;
        352 : storage = 256'h583e25abe62029417f47229b4c634219876e48be79199e7d070dcf9a0d49ef61;
        353 : storage = 256'h0e7449695d6309a0d28b83a87e0ea881104e393d282be26894b6aa57a9d312bf;
        354 : storage = 256'h11090e110867b17b19f13a7184638de12d4429c9ed7d91ed53c2d2e8e2dd0e11;
        355 : storage = 256'h15dcf29ad129c47d27414803871eefb91e8f377758f374e67865daa06e054137;
        356 : storage = 256'h040bc6cc790bb5180a8010b4af71dea5866550de1d58e5e49773e7e30122f1a1;
        357 : storage = 256'h281792399e8ca15cedee0277f5c22b81739777e06274e0ae25957e26b249521b;
        358 : storage = 256'h32416530c61380069621c68f25024ba56e2298b83fa864b19d371a6f592ee1f9;
        359 : storage = 256'h0bf30c2917230163e3b6348def8c8fbd0c28d06cf4a8ff26edc26e72c42cc665;
        360 : storage = 256'h74081ee0cfa7f006498ccd02b132f0317d608896cb6977d16ce452622cc0fd79;
        361 : storage = 256'h2ee2823585f35456ad45f5dcfff449f57aec1ccc75209f0d40d311d21128a939;
        362 : storage = 256'h2851e9388b3003a7524ec53f5e838d213137f7cf6c2f865a217121d0c0763c4d;
        363 : storage = 256'h66b5525f39a54f9ea8684f07e1eb674970b5ed8b53d173f63d3f85a2e8a32f77;
        364 : storage = 256'h2d5a4e381a5033aa87004d4f3fac178175a02d3fc7acbe4aff7d80167a20729b;
        365 : storage = 256'h534e0f35bc56936607d9962f6a2ff1499ec954cbb4e4473fe6a46b4dd6b0999f;
        366 : storage = 256'h699ab1c1acf857cdb4f7b00074d57b6980e0ad6d4d65db4078e1cd847cc96f2d;
        367 : storage = 256'h010d66408231f6391d8ad93cd8f9464102ccc6b12f2b12a8bbb5cf65b884f13f;
        368 : storage = 256'h650119f1c9764b2f807a2bdfb460f4656bfdac6d04971673cc3048a93df03bd9;
        369 : storage = 256'h7179a3110af4eb0d834287d22e274bf1857236f17ac3edc552dc71307ad630a3;
        370 : storage = 256'h6bb5ab655bf358c623e2ac325173071d9fd6c4c4f7e4fdd74ee6ae5343303c91;
        371 : storage = 256'h06e187c413614ebca34dba6666d59f9919e083b412002d920c2f36f5703dd777;
        372 : storage = 256'h111daef262d51b7e957669cbc6e68e5971513b4d30a1be9182c45edd2f229a9f;
        373 : storage = 256'h4fedd9d326dfa2236f69a8fa655f9ff16238102bdb3ec173845ff52a276c55fb;
        374 : storage = 256'h0d67d4fc9bd3044e63e9698239a1039d17079e7c4c4185c2a51b7602f702e705;
        375 : storage = 256'h009608f7ac043eef37784dbbbfda67a108c90cbf69dc925b8e79229d2499683f;
        376 : storage = 256'h22b8325b9c5321bc579c89d1e97c9a49572243497dc329819221ccd14c94d6b9;
        377 : storage = 256'h9a3a21aa91a68b132aadcbd7dd75a809b601ce79c4deea100f17ee78eb78d38d;
        378 : storage = 256'h1ac5a49edf23422595c88fcac0b21eb14023549a1b5876f8df7477a2c69a13d1;
        379 : storage = 256'h0a6e0b6fd0ee65cb3b48731ddddc6ddd0e39d6c2e830d6e0095ecd8409ff3dcd;
        380 : storage = 256'h10ebcae521abf6f5a3ca08b9f15d3781189987e32d7b64757e6d01c44ca825ab;
        381 : storage = 256'h56fc96358cf85dd41ff23f1b6dd708b19cad4870b4a9537eb096286793526d97;
        382 : storage = 256'h0265d76e68e11a152aa1c2d57f0d7c611630812131f058b85bca878560ab2edb;
        383 : storage = 256'h583e25abe62029417f47229b4c634219876e48be79199e7d070dcf9a0d49ef61;
        384 : storage = 256'h06006058320c617cd4fc6a3fe991bc611041692c813655d7d4ab5fb1fa6ff877;
        385 : storage = 256'h17ad6c489e11c7011422717d084933092d2097ebb53629820ac41d59029762d9;
        386 : storage = 256'h0e7ffdaedb6cca9d2fb7540d12f847c11e77340ea69a9bb1ca9f80c693ec38af;
        387 : storage = 256'h316b4765e47e69cdd9a324401f76f2f585fbb57fb5269adc374a8184125b46e9;
        388 : storage = 256'h3d5708b1de5061b88e0df07735e84a81733ca32ee837d4aface667f7dfca89b3;
        389 : storage = 256'h316f351cfc341b69da7e99feb46a157d6dcc0dacc6573969ccca429d14a3d001;
        390 : storage = 256'h01c5b841d59bff4072a13c073f4637090c1f4267ecb4bc3534e056a1d51272cd;
        391 : storage = 256'h031dca3429c0324f2b70d11bd6d12f297cfe03707b834cacc1d533fc2f9da781;
        392 : storage = 256'h383633bb86b9c8315eb0a1e60c860c197a8b8574ce4320fcf6f753bd9f95a141;
        393 : storage = 256'h0417a7210f45cd7fbf6d7db6f7b27f3931114ae02bc8c5586d78f16c877c11f5;
        394 : storage = 256'h4a7b0811fd314d6512fae92ad6267469705d5c6734dfc942cf7d830aa64d28ef;
        395 : storage = 256'h19a30e1cb2be17205ea8e4dd2d3ee4017543bf635b3e5a998b93d1796c52ce33;
        396 : storage = 256'h3e8053dfb582d342d70c199203a2fae19e4c8ef0761ca8a509d8b3b2572f6e57;
        397 : storage = 256'h4f099b93e22ba71ffe40d68aa1a47ed1807b681892801f5f194dff894d4993d5;
        398 : storage = 256'h0010cd58d0c69dea39a972d0d13e337902ca9374ce90f9ff027aa68e32986af7;
        399 : storage = 256'h0a4385e2899126b24a444d0f0ce288216ba8d0b83151a116a69a638c287a70e1;
        400 : storage = 256'h76b2f3dda02fa9cb31bcaf3c494051e185095a99e56c1e8f25b67aea35a8fe7b;
        401 : storage = 256'h45f7792789a91de31990647023019ca19f592b310fbc073b5e6bcfdb7fbfa559;
        402 : storage = 256'h058417fa1556e48906888b4fa2f3074919cc2e3921d5526987253098906710ef;
        403 : storage = 256'h00dbc77b1bb65ee1124de383f96b81410da4a54cec79d4444f08b9940aada341;
        404 : storage = 256'h0166207f2ce2dcdd9a9f7801aa37ec210bd349c68696b155187f56839aaa3b65;
        405 : storage = 256'h01ee62275c4c59d0ece4a1a274eab67102c5d1b4ff0005e8726d78b245cc279b;
        406 : storage = 256'h00b8660d19ae53911bbac1d2d0aacd21010ec7ce87df4fc9280567c6f27449a1;
        407 : storage = 256'h014dc59551fb9b9b3b6ec0938be815d90a7d9f9b286ac98f505a59fcd4a8a667;
        408 : storage = 256'h048fb7d0fc9499327f96dd3b8a7f099115e9c9e4af4cdc11e527eeec97ed7c13;
        409 : storage = 256'h05f534d603e3d9a902360d97a90ed2e107b8d9a3bcd094256e6ebbc726bd1c4f;
        410 : storage = 256'h0079094049ca53307b452d0f8161aab901b67819f7932ab464bfe21c6005d9d3;
        411 : storage = 256'h013d89f5322b7d74d76a0869a372252102f6355b90a42723ec2cc968274581b5;
        412 : storage = 256'h10c05e85391d1dcb0572fbbbdbc3af7112dd11140f94e9c95186e790e0b37f49;
        413 : storage = 256'h01f503baf4c64d09296e422133586a4102abeb7b406e3cc3923cfe186e11be85;
        414 : storage = 256'h0e7449695d6309a0d28b83a87e0ea881104e393d282be26894b6aa57a9d312bf;
        415 : storage = 256'h06006058320c617cd4fc6a3fe991bc611041692c813655d7d4ab5fb1fa6ff877;
        416 : storage = 256'h0379ad6405d469677492f48e4bd4aa01056ee7f306350d43bcd7dd94789a5e47;
        417 : storage = 256'h01fce5d04c5bc615540227155196b52103ab01a335dec6adf848814065792731;
        418 : storage = 256'h05c11743877cbe02a9a304b3d469e1b110219b700dab4db919c08a9856385c37;
        419 : storage = 256'h060970482c38138a1b47e933f2cfac010ddfcf522a728cb767b216479a2e4ead;
        420 : storage = 256'h0066236a6e8c7505ae444723282d93310d38255909f38511693b384c99fb061f;
        421 : storage = 256'h006d7e3bd3dbc2f4a095862564c530f10175a019d549b1ca4bf22e0619a744d3;
        422 : storage = 256'h027791a63d042890b6f45dafd1a92c410f0c7cfe40ad36d39263fbb5f6611e9f;
        423 : storage = 256'h0b29c3a894578c74c2b6f727cba9d9710ec10f5db97a3f672e798b63a72edcdf;
        424 : storage = 256'h052082aaab86756d7e454df97192622905e859e39be2db301e553a8ed61cfaab;
        425 : storage = 256'h09166f925622ca6d84723e3e10c37c810d8748c30b9d0230e14d24b5f90bbef1;
        426 : storage = 256'h02b41f2c8c2c5eb3a0382a20d9b8de010e1e4f3db656f4b3b66c4440b9f19a2d;
        427 : storage = 256'h033253a75a60b9dd92005748d81c9f01130f109f11b3b56fe344983d0a171689;
        428 : storage = 256'h036bac9410bcbf0e24ff8a0863586fe10f780cff2ce21b7855ec1871d410f4cb;
        429 : storage = 256'h000a246b5da499317bfab9bbba6b0be10056088851a4a4492ba9be53b97b6de9;
        430 : storage = 256'h0b403160b96fb4eda5f20c05bd38c0590cf64279428c49058da419a4e6f3c13f;
        431 : storage = 256'h01558d17df1fdb72e4285d63b438916110046d9d0fca79070587cfcdcadda2e5;
        432 : storage = 256'h073ffcd060e991ecd8851f54ee6a4851132f67ae70b0d4434a59107bf2116bc7;
        433 : storage = 256'h0169aea9f0fea53f357eebcdd354da51031b20dc628def68a14877889a1ed6f1;
        434 : storage = 256'h1d324b6d3b6a9ca0f6b978455a50d8c125e004b336e3615048b21910b6a65bef;
        435 : storage = 256'h1c57c8eef87f7abad3a1748cf377922120d420c98aaa832abdb6a3641591368b;
        436 : storage = 256'h01f42d0faf9e2f6b872d01d44a49ee8507b28bd312e9511d1b8433f0da33f675;
        437 : storage = 256'h00dcd8b9ac6da812c32fd7d022b07fb102efb8651e1ea3f8e33a5d7a992e078f;
        438 : storage = 256'h0a04c4065adecaca84179fcc88f275851d1f9fd5d662a6246bf976b4d28f21e9;
        439 : storage = 256'h00c4c1ac8b5e2f04171eab9c4d6027113cd5785d1364e935d2f76f73cc02e07d;
        440 : storage = 256'h030654df9a1b6b7686c3d8026568a02d156ffb4ab15220e3e2926b27cb9b7f81;
        441 : storage = 256'h03ec0a706df78f5cd5b566e2b8a2e05904c13eac83289c1bf62ba243016d56bd;
        442 : storage = 256'h014384dca78c888a239b60f7318898510838e17b4bca6db519e1d9853bc80f3b;
        443 : storage = 256'h1e0fdd5c1c59ff328605373eb15c6c11345e16cf01638c15f85585f1b16ad967;
        444 : storage = 256'h055e4eb8a2292817324478e463dc8121076aa57ea3b2637e571f857f096fa96b;
        445 : storage = 256'h11090e110867b17b19f13a7184638de12d4429c9ed7d91ed53c2d2e8e2dd0e11;
        446 : storage = 256'h17ad6c489e11c7011422717d084933092d2097ebb53629820ac41d59029762d9;
        447 : storage = 256'h0379ad6405d469677492f48e4bd4aa01056ee7f306350d43bcd7dd94789a5e47;
        448 : storage = 256'h059949a486cd30c2134d27ef42f797510a2ecc646e544fd98f668bce81d564ff;
        449 : storage = 256'h0a9172859be413e7a53df04e429a9f692cc84d73254559f1f3e92d3edb24f319;
        450 : storage = 256'h14a3c5ffb8019bb517cc8994b516ab81268443ef3838119af7610e70256f98c3;
        451 : storage = 256'h0a5d6e647431e1e26838f9154851935924b2cf3473ee45450bcfba84fa48dcb1;
        452 : storage = 256'h007d0bd9341f621c247a26098367950d040d3b029fa04b8b7d34ecb4ce30fbbd;
        453 : storage = 256'h13302efcc957555c8294683b1856788529c6fc6927a88f870f272f2fc420dc31;
        454 : storage = 256'h0f2cff36f4291823d92030391ff045c928f5967cbc563e4211d5724858c989f1;
        455 : storage = 256'h0af20966f2e347b8dac71b48eea0d3e51066798011aa572d055916efb99de665;
        456 : storage = 256'h1a0cb3733757cf10e7962e3d4c9d38a9258e81daece5bde144ac0697339e813f;
        457 : storage = 256'h1a67b5c16959838530fa0a992a8ac4012731c5b3460f02bb8dbc9acaeddcf543;
        458 : storage = 256'h2ff2de9ce65c2590a7d1bdd56354c00134e8e3ee172477180c66a89cedc15e27;
        459 : storage = 256'h087d7d5177acec60061d95715dca16fd2af197c709dde63807225634c20b3245;
        460 : storage = 256'h000aa349059860c0e856ccf880f00de900eed6d698325f01ab496c7a00ef88c7;
        461 : storage = 256'h0e165b1ab32714137b02466a960a7f1523fbe6aabe0dfb2df64ffc11de789791;
        462 : storage = 256'h154ea533fa776cd2565fa34050a096412c774c4a3627e7d2cffa139a5867b70b;
        463 : storage = 256'h138435be15a9ca95b57822c83466a83d3542aba113b582b3870ebab714977e89;
        464 : storage = 256'h0560c25850dfc87b4ce3e3fd6a3daae1089f600755cd344d92c87a1cb667e93f;
        465 : storage = 256'h0ee51c5c9eda7e51c74bc9150785d7d11991d2666a8bd1dec96ac95ff1d624c9;
        466 : storage = 256'h111080f4f29036718f3e9d5d54193f611629a95384a003bededde0953d588c0d;
        467 : storage = 256'h03198ab43d875dbdc9ef49f87e8ebcd9053252e704e0448ee9630f4957b76ef3;
        468 : storage = 256'h00b1381299ba2bbef467e586497081e101fb7d4d5bfa9a3e8a606bc09ed1ce29;
        469 : storage = 256'h00e9efc2e9b343a0bcd8090feab381f113a9529a6dc6f615d9f8a5d337d2de1f;
        470 : storage = 256'h0c9886363201a143c4306bf30986c1612911b6b9718e06b2323a288a1cc4eb2b;
        471 : storage = 256'h0c06a3283717e2ea451e9534ca6ee3510e78f57e2c2b7bac583a24022d374f47;
        472 : storage = 256'h01efaa713b6b315ce2cfada561e814710335c45918e247a0865c44cf299f56eb;
        473 : storage = 256'h01ce45fd539233703f24c997c6ce7901058d03805addfb9c9deb7a73754d5cdd;
        474 : storage = 256'h1d7c243ac2b170d82fa472a8b73cd5e1235a8181f77ed27ee31ec51e25951d11;
        475 : storage = 256'h03e070bef1c25eb620c72ac3e9d7cda10501c8b6a48b969a535bcbe483b3982d;
        476 : storage = 256'h15dcf29ad129c47d27414803871eefb91e8f377758f374e67865daa06e054137;
        477 : storage = 256'h0e7ffdaedb6cca9d2fb7540d12f847c11e77340ea69a9bb1ca9f80c693ec38af;
        478 : storage = 256'h01fce5d04c5bc615540227155196b52103ab01a335dec6adf848814065792731;
        479 : storage = 256'h059949a486cd30c2134d27ef42f797510a2ecc646e544fd98f668bce81d564ff;
        480 : storage = 256'h17c8a0e302be3793f2cf8e2dd586bb091e3b99093fa8436c972a745cac23da6f;
        481 : storage = 256'h051d906d1d2d13b485557f9fd94579011a00b4a933e30733e4a59553fae5d595;
        482 : storage = 256'h03fa7b2ec67c0c0c1fb59ee2c4512ce118c6797674d491601a9a176c172e1f97;
        483 : storage = 256'h005aab75f16feea54765e5bdac4c2d1102bc3d13c1aba79638edac9bbbee99eb;
        484 : storage = 256'h015bcebb38e4e2f75939f84b637ee7a91c343aa156880e9e53f09ebaf5fcbc17;
        485 : storage = 256'h0f7832826b2baa02170a4c9c141e69c11ba6dd0cffb512ec71238a7b7b0b4c57;
        486 : storage = 256'h03fe3b88ec551c19ad6e4f8a1fa0d4610b1268507e7be91d14d502f8acedd283;
        487 : storage = 256'h03f75c06739592e7b36cff87ac9f9ec1195acb1b7543621eb103fbbfe104c5f9;
        488 : storage = 256'h02da703364e492e369e458ef31eb49011a75d74700fa1663b7619b439bf9bd15;
        489 : storage = 256'h03987670be7bac92f37567afe13b2fb123b83610696979c2d9a447ed06c3ce51;
        490 : storage = 256'h14a75ab7f61f62370d0a52e803c278391cfdd1dc8d0b1db7f56b6940c4b58da3;
        491 : storage = 256'h006138bb58ce82e4c587305a9bdb544100a13dc816a9158119fefe7099fa30b1;
        492 : storage = 256'h00f74a6e99980f9e5d3628793ffeda71184afe064a224e0b0a7a3ecc8cc823b7;
        493 : storage = 256'h0889db15c9d63c7cf9e4681993fd82e11e04e94b4fc6bcb6bd42a5094f2f6f8d;
        494 : storage = 256'h040d856739ecb943edfa55f59f35a5b923f4d274360f91210d12cd5ab46a1e7f;
        495 : storage = 256'h02edaf90a448b481f861e5d64875c5a105d235409db9c86567b3923161e49df9;
        496 : storage = 256'h2d1f8eadbf09df92173771be025fa1d17073872fe431bfe990e5ef77fd90185f;
        497 : storage = 256'h53e12b6aa2acc70fafd8bd0c07aeef016177e6330bcc7b28c9b0ad3fb200c2bb;
        498 : storage = 256'h13822f0e1b7a0515476382890c7b316116da8fcc36121641fd9f1280fa7fba45;
        499 : storage = 256'h088897d3de8f3417e8a880509a1eaf6908b7dc8436b787004bc8f07f983e8dff;
        500 : storage = 256'h527dc71a041c8b0216f63ea699a72fcd5677c96d81061c07aaae244cae9a1ef9;
        501 : storage = 256'h35b31251dea063a0723f6b10c51000adb49db6695afc781a0e73035800d918cd;
        502 : storage = 256'h25af78db5925d4ae5cbcfb764c658e113fa5d86f5ffc14827ca18977ef229211;
        503 : storage = 256'h0132298fa9c1c9a8f74abd9812868f410e1e018f46e41f7c0bb2fffe26b8930d;
        504 : storage = 256'h086d5a756222e70d85bb7cb787ca9e01186966dd90069f25ee621cfab87f5e6b;
        505 : storage = 256'h889c0653bf0caf00a68ecc6494401aa99b7abf3f1d172ac698eea2c28b175957;
        506 : storage = 256'h117f422294915e573434e6ee19c533411605174f7440323a12d336ce13e2939b;
        507 : storage = 256'h040bc6cc790bb5180a8010b4af71dea5866550de1d58e5e49773e7e30122f1a1;
        508 : storage = 256'h316b4765e47e69cdd9a324401f76f2f585fbb57fb5269adc374a8184125b46e9;
        509 : storage = 256'h05c11743877cbe02a9a304b3d469e1b110219b700dab4db919c08a9856385c37;
        510 : storage = 256'h0a9172859be413e7a53df04e429a9f692cc84d73254559f1f3e92d3edb24f319;
        511 : storage = 256'h17c8a0e302be3793f2cf8e2dd586bb091e3b99093fa8436c972a745cac23da6f;
    endcase
    
    case (storage3)
        0 : p3 = 32'd17627;
        1 : p3 = 32'd32423;
        2 : p3 = 32'd63863;
        3 : p3 = 32'd51853;
        4 : p3 = 32'd36571;
        5 : p3 = 32'd38501;
        6 : p3 = 32'd60271;
        7 : p3 = 32'd25097;
        8 : p3 = 32'd62081;
        9 : p3 = 32'd31397;
        10 :p3 = 32'd49339;
        11 :p3 = 32'd19507;
        12 :p3 = 32'd22129;
        13 :p3 = 32'd43177;
        14 :p3 = 32'd11833;
        15 :p3 = 32'd26813;
        16 :p3 = 32'd3137;
        17 :p3 = 32'd27259;
        18 :p3 = 32'd60343;
        19 :p3 = 32'd751;
        20 :p3 = 32'd58453;
        21 :p3 = 32'd56873;
        22 :p3 = 32'd22307;
        23 :p3 = 32'd28901;
        24 :p3 = 32'd14897;
        25 :p3 = 32'd30013;
        26 :p3 = 32'd52433;
        27 :p3 = 32'd56197;
        28 :p3 = 32'd7331;
        29 :p3 = 32'd25759;
        30 :p3 = 32'd13477;
        31 :p3 = 32'd25243;
    endcase
    
    case (storage4)
        0 : p4 = 32'd17627;
        1 : p4 = 32'd32423;
        2 : p4 = 32'd63863;
        3 : p4 = 32'd51853;
        4 : p4 = 32'd36571;
        5 : p4 = 32'd38501;
        6 : p4 = 32'd60271;
        7 : p4 = 32'd25097;
        8 : p4 = 32'd62081;
        9 : p4 = 32'd31397;
        10 :p4 = 32'd49339;
        11 :p4 = 32'd19507;
        12 :p4 = 32'd22129;
        13 :p4 = 32'd43177;
        14 :p4 = 32'd11833;
        15 :p4 = 32'd26813;
        16 :p4 = 32'd3137;
        17 :p4 = 32'd27259;
        18 :p4 = 32'd60343;
        19 :p4 = 32'd751;
        20 :p4 = 32'd58453;
        21 :p4 = 32'd56873;
        22 :p4 = 32'd22307;
        23 :p4 = 32'd28901;
        24 :p4 = 32'd14897;
        25 :p4 = 32'd30013;
        26 :p4 = 32'd52433;
        27 :p4 = 32'd56197;
        28 :p4 = 32'd7331;
        29 :p4 = 32'd25759;
        30 :p4 = 32'd13477;
        31 :p4 = 32'd25243;
    endcase
end

endmodule            